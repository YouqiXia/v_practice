package dut_package;
    typedef struct{
        int addr;
        int data;
    }tx_packet_t;

endpackage